module sky130_fd_sc_hd__bufbuf_16 (
    X,
    A
);

    output X   ;
    input  A   ;

    assign X = A;
endmodule
